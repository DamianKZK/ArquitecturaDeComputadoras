module adder(
	input [32:0]pcIn,
	output [32:0]pcOut);
	
	assign pcOut = pcIn+4;

endmodule