`timescale 1ns/1ns
module shiftLeft2(
	input inData,
	output outData);

assign outData = inData<<2;


endmodule