//1.Definición del modulo y sus entradas y salidas
//https://github.com/DamianKZK/ArquitecturaDeComputadoras/upload

module _and(input A, input B, output C);
//2. Declarar señales/elementos internos

//3.Comportamiento del modulo (asignaciones, instancias y conexiones)

assign C=A&B;
endmodule